module not_gate(x,y);
input x;
output y;
assign y = ~x;
endmodule